package i2c_agent_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  
  `include "i2c_sequence_item.sv"
endpackage
