package i2c_agent_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "defines.sv"
  `include "i2c_sequence_item.sv"
  `include "i2c_agent_config.sv"
  `include "i2c_monitor.sv"  
  `include "i2c_agent.sv"  
endpackage