package wb_i2c_seq_pkg;
  import uvm_pkg::*;

  `include "wb_i2c_seq.sv"
endpackage