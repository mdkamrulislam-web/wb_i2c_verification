// ########################### \\
// Register Address Definition \\
// ########################### \\

`define PRER_LO 3'b000
`define PRER_HI 3'b001
`define CTR     3'b010
`define TXR     3'b011
`define CR      3'b100
`define RXR     3'b011
`define SR      3'b100
`define SLVADDR 7'h3C 
`define WR      1'b0  
`define RD      1'b1  