package wb_agent_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"
  
  `include "defines.sv"
  `include "wb_sequence_item.sv"
  `include "wb_agent_config.sv"
  `include "wb_driver.sv"
  `include "wb_monitor.sv"
  `include "wb_sequencer.sv"

  `include "wb_agent.sv"
  
endpackage